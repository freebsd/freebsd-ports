share/aspell/sv.dat
share/aspell/sv.multi
share/aspell/sv.rws
share/aspell/sv_phonet.dat
share/aspell/svenska.alias
share/aspell/swedish.alias
