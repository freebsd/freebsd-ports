lib/aspell-%%VER%%/sv_phonet.dat
lib/aspell-%%VER%%/sv.dat
share/aspell/sv.multi
share/aspell/sv.rws
share/aspell/svenska.alias
share/aspell/swedish.alias
