usr/lib/aspell/sv.multi
usr/lib/aspell/sv.rws
usr/lib/aspell/svenska.alias
usr/lib/aspell/swedish.alias
usr/share/aspell/sv.dat
usr/share/aspell/sv_phonet.dat
